module hash_round (
   
);
   
	// Declarations
	
	// State splitting
	
	// Mix function
	
	// Rotator
	
	// Output state assignment

endmodule
