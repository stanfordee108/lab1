module hash_rom(
   
);
   
	// Module body

endmodule
