module cam (
      
);
	// wire declarations

	// data concatenation
	
	// 8 equality comparisons
	
	// encoder instantiation
	
	// valid logic
	
endmodule
