module arbiter (
   
);
   
	// module body goes here

endmodule
