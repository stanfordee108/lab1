module hasher (
   
);

	// DO IT GORDON
	
endmodule
