module verifier (
   
);

	// FINISH HIM

endmodule
