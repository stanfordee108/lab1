module length_finder (
   
);
   
	// wire declarations
	
	// is_character_null logic (8 lines of it!)
	
	// arbiter
  
endmodule
