module encoder (
   
);
   
endmodule
